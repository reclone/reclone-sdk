//
// 6502DecodeRom - ROM acting as a lookup table to decode 6502 opcodes into CPU control signals.
//
//
// Copyright 2018 Reclone Labs <reclonelabs.com>
// 
// Redistribution and use in source and binary forms, with or without modification, are permitted
// provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this list of
//    conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice, this list of
//    conditions and the following disclaimer in the documentation and/or other materials
//    provided with the distribution.
// 
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR
// IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND
// FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
// CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR 
// OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.

module Cpu6502DecodeRom
(
    input                       clock,
    input                       enable,
    input [7:0]                 address,
    output reg [31:0]           data
);

parameter CYC0_INCREMENT_PC         =   32'h00000001;
parameter CYC1_INCREMENT_PC         =   32'h00000002;

parameter ALU_OPERAND1_IS_ZERO      =   32'h00000000;
parameter ALU_OPERAND1_IS_A         =   32'h00000004;
parameter ALU_OPERAND1_IS_X         =   32'h00000008;
parameter ALU_OPERAND1_IS_Y         =   32'h0000000C;

parameter ALU_OPERAND2_IS_ZERO      =   32'h00000000;
parameter ALU_OPERAND2_IS_IMM       =   32'h00000010;

parameter ALU_OPERATION_IS_ASSIGN   =   32'h00000000;

parameter STORE_ALU_OUTPUT_NOWHERE  =   32'h00000000;
parameter STORE_ALU_OUTPUT_IN_A     =   32'h00001000;

always @ (posedge clock)
begin
    if (enable)
    begin
        case (address)
            8'hA9:   //LDA #immediate
                data <= CYC0_INCREMENT_PC;
            default: //NOP
                data <= 0;
        endcase
    end
end


endmodule
